// HPS.v

// Generated using ACDS version 14.0 200 at 2018.12.24.16:01:26

`timescale 1 ps / 1 ps
module HPS (
		output wire [14:0] memory_mem_a,                     // memory.mem_a
		output wire [2:0]  memory_mem_ba,                    //       .mem_ba
		output wire        memory_mem_ck,                    //       .mem_ck
		output wire        memory_mem_ck_n,                  //       .mem_ck_n
		output wire        memory_mem_cke,                   //       .mem_cke
		output wire        memory_mem_cs_n,                  //       .mem_cs_n
		output wire        memory_mem_ras_n,                 //       .mem_ras_n
		output wire        memory_mem_cas_n,                 //       .mem_cas_n
		output wire        memory_mem_we_n,                  //       .mem_we_n
		output wire        memory_mem_reset_n,               //       .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                    //       .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                   //       .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                 //       .mem_dqs_n
		output wire        memory_mem_odt,                   //       .mem_odt
		output wire [3:0]  memory_mem_dm,                    //       .mem_dm
		input  wire        memory_oct_rzqin,                 //       .oct_rzqin
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO01, // hps_io.hps_io_gpio_inst_LOANIO01
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO02, //       .hps_io_gpio_inst_LOANIO02
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO03, //       .hps_io_gpio_inst_LOANIO03
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO04, //       .hps_io_gpio_inst_LOANIO04
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO05, //       .hps_io_gpio_inst_LOANIO05
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO06, //       .hps_io_gpio_inst_LOANIO06
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO07, //       .hps_io_gpio_inst_LOANIO07
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO08, //       .hps_io_gpio_inst_LOANIO08
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO10, //       .hps_io_gpio_inst_LOANIO10
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO11, //       .hps_io_gpio_inst_LOANIO11
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO12, //       .hps_io_gpio_inst_LOANIO12
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO13, //       .hps_io_gpio_inst_LOANIO13
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO42, //       .hps_io_gpio_inst_LOANIO42
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO49, //       .hps_io_gpio_inst_LOANIO49
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO50, //       .hps_io_gpio_inst_LOANIO50
		output wire [66:0] loanio_in,                        // loanio.in
		input  wire [66:0] loanio_out,                       //       .out
		input  wire [66:0] loanio_oe,                        //       .oe
		input  wire [31:0] hps_gp_gp_in,                     // hps_gp.gp_in
		output wire [31:0] hps_gp_gp_out                     //       .gp_out
	);

	HPS_hps_0 #(
		.F2S_Width (0),
		.S2F_Width (0)
	) hps_0 (
		.h2f_loan_in               (loanio_in),                        // h2f_loan_io.in
		.h2f_loan_out              (loanio_out),                       //            .out
		.h2f_loan_oe               (loanio_oe),                        //            .oe
		.h2f_gp_in                 (hps_gp_gp_in),                     //      h2f_gp.gp_in
		.h2f_gp_out                (hps_gp_gp_out),                    //            .gp_out
		.mem_a                     (memory_mem_a),                     //      memory.mem_a
		.mem_ba                    (memory_mem_ba),                    //            .mem_ba
		.mem_ck                    (memory_mem_ck),                    //            .mem_ck
		.mem_ck_n                  (memory_mem_ck_n),                  //            .mem_ck_n
		.mem_cke                   (memory_mem_cke),                   //            .mem_cke
		.mem_cs_n                  (memory_mem_cs_n),                  //            .mem_cs_n
		.mem_ras_n                 (memory_mem_ras_n),                 //            .mem_ras_n
		.mem_cas_n                 (memory_mem_cas_n),                 //            .mem_cas_n
		.mem_we_n                  (memory_mem_we_n),                  //            .mem_we_n
		.mem_reset_n               (memory_mem_reset_n),               //            .mem_reset_n
		.mem_dq                    (memory_mem_dq),                    //            .mem_dq
		.mem_dqs                   (memory_mem_dqs),                   //            .mem_dqs
		.mem_dqs_n                 (memory_mem_dqs_n),                 //            .mem_dqs_n
		.mem_odt                   (memory_mem_odt),                   //            .mem_odt
		.mem_dm                    (memory_mem_dm),                    //            .mem_dm
		.oct_rzqin                 (memory_oct_rzqin),                 //            .oct_rzqin
		.hps_io_gpio_inst_LOANIO01 (hps_io_hps_io_gpio_inst_LOANIO01), //      hps_io.hps_io_gpio_inst_LOANIO01
		.hps_io_gpio_inst_LOANIO02 (hps_io_hps_io_gpio_inst_LOANIO02), //            .hps_io_gpio_inst_LOANIO02
		.hps_io_gpio_inst_LOANIO03 (hps_io_hps_io_gpio_inst_LOANIO03), //            .hps_io_gpio_inst_LOANIO03
		.hps_io_gpio_inst_LOANIO04 (hps_io_hps_io_gpio_inst_LOANIO04), //            .hps_io_gpio_inst_LOANIO04
		.hps_io_gpio_inst_LOANIO05 (hps_io_hps_io_gpio_inst_LOANIO05), //            .hps_io_gpio_inst_LOANIO05
		.hps_io_gpio_inst_LOANIO06 (hps_io_hps_io_gpio_inst_LOANIO06), //            .hps_io_gpio_inst_LOANIO06
		.hps_io_gpio_inst_LOANIO07 (hps_io_hps_io_gpio_inst_LOANIO07), //            .hps_io_gpio_inst_LOANIO07
		.hps_io_gpio_inst_LOANIO08 (hps_io_hps_io_gpio_inst_LOANIO08), //            .hps_io_gpio_inst_LOANIO08
		.hps_io_gpio_inst_LOANIO10 (hps_io_hps_io_gpio_inst_LOANIO10), //            .hps_io_gpio_inst_LOANIO10
		.hps_io_gpio_inst_LOANIO11 (hps_io_hps_io_gpio_inst_LOANIO11), //            .hps_io_gpio_inst_LOANIO11
		.hps_io_gpio_inst_LOANIO12 (hps_io_hps_io_gpio_inst_LOANIO12), //            .hps_io_gpio_inst_LOANIO12
		.hps_io_gpio_inst_LOANIO13 (hps_io_hps_io_gpio_inst_LOANIO13), //            .hps_io_gpio_inst_LOANIO13
		.hps_io_gpio_inst_LOANIO42 (hps_io_hps_io_gpio_inst_LOANIO42), //            .hps_io_gpio_inst_LOANIO42
		.hps_io_gpio_inst_LOANIO49 (hps_io_hps_io_gpio_inst_LOANIO49), //            .hps_io_gpio_inst_LOANIO49
		.hps_io_gpio_inst_LOANIO50 (hps_io_hps_io_gpio_inst_LOANIO50), //            .hps_io_gpio_inst_LOANIO50
		.h2f_rst_n                 ()                                  //   h2f_reset.reset_n
	);

endmodule
