// asmi.v

// Generated using ACDS version 14.0 200 at 2018.10.27.20:17:39

`timescale 1 ps / 1 ps
module asmi (
		input  wire        clkin,      //      clkin.clk
		input  wire        read,       //       read.read
		input  wire        rden,       //       rden.rden
		input  wire [23:0] addr,       //       addr.addr
		input  wire        reset,      //      reset.reset
		output wire [7:0]  dataout,    //    dataout.dataout
		output wire        busy,       //       busy.busy
		output wire        data_valid  // data_valid.data_valid
	);

	asmi_asmi_parallel_0 asmi_parallel_0 (
		.clkin      (clkin),      //      clkin.clk
		.read       (read),       //       read.read
		.rden       (rden),       //       rden.rden
		.addr       (addr),       //       addr.addr
		.reset      (reset),      //      reset.reset
		.dataout    (dataout),    //    dataout.dataout
		.busy       (busy),       //       busy.busy
		.data_valid (data_valid)  // data_valid.data_valid
	);

endmodule
