
module clock_control (
	inclk,
	ena,
	outclk);	

	input		inclk;
	input		ena;
	output		outclk;
endmodule
